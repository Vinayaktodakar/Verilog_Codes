module ripple_carry_adder_4bit (
    input  [3:0] A,    // 4-bit input operand A
    input  [3:0] B,    // 4-bit input operand B
    input        cin,  // Initial carry-in (usually 0)
    output [3:0] Sum,  // 4-bit result sum
    output       cout  // Final carry-out
);
    // Intermediate carry signals
    wire c1, c2, c3;

    // Instantiate 4 Full Adders
    full_adder FA0 (.a(A[0]), .b(B[0]), .cin(cin), .sum(Sum[0]), .cout(c1));
    full_adder FA1 (.a(A[1]), .b(B[1]), .cin(c1),  .sum(Sum[1]), .cout(c2));
    full_adder FA2 (.a(A[2]), .b(B[2]), .cin(c2),  .sum(Sum[2]), .cout(c3));
    full_adder FA3 (.a(A[3]), .b(B[3]), .cin(c3),  .sum(Sum[3]), .cout(cout));

endmodule
